// Build ID Verilog Module
`define BUILD_DATE "20230427"
`define BUILD_HASH "a36b0dad"
